
package bp_be_hardfloat_pkg;

localparam dword_width_gp  = 64;
localparam word_width_gp   = 32;

localparam float_width_gp  = 32;
localparam double_width_gp = 64;



endpackage

